/********************************************************************************************

Filename:	async_fifo_package.sv   

Description:	package for async fifo testbench 

Version:	1.0

*********************************************************************************************/


package fifo_pkg;

`include "seq_item.sv"
`include "seq_base.sv"
`include "seq_full.sv"
`include "seq_random.sv"

`include "sequencer.sv"
`include "driver.sv"
`include "write_monitor.sv"
`include "read_monitor.sv"
`include "write_agent.sv"
`include "read_agent.sv"
`include "scoreboard.sv"

		
endpackage:fifo_pkg

